-- audioInTest.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity audioInTest is
	port (
		reg_clk     : in  std_logic                     := '0';             --       control_clock.clk
		reg_reset   : in  std_logic                     := '0';             -- control_clock_reset.reset
		aes_clk     : in  std_logic                     := '0';             --   conduit_aes_audio.export
		aes_de      : in  std_logic                     := '0';             --                    .export
		aes_ws      : in  std_logic                     := '0';             --                    .export
		aes_data    : in  std_logic                     := '0';             --                    .export
		aud_clk     : in  std_logic                     := '0';             --          dout_clock.clk
		reset       : in  std_logic                     := '0';             --    dout_clock_reset.reset
		aud_ready   : in  std_logic                     := '0';             --                dout.ready
		aud_valid   : out std_logic;                                        --                    .valid
		aud_sop     : out std_logic;                                        --                    .startofpacket
		aud_eop     : out std_logic;                                        --                    .endofpacket
		aud_channel : out std_logic_vector(7 downto 0);                     --                    .channel
		aud_data    : out std_logic_vector(23 downto 0);                    --                    .data
		channel0    : in  std_logic_vector(7 downto 0)  := (others => '0'); --     conduit_control.export
		channel1    : in  std_logic_vector(7 downto 0)  := (others => '0'); --                    .export
		fifo_status : out std_logic_vector(7 downto 0);                     --                    .export
		fifo_reset  : in  std_logic                     := '0'              --                    .export
	);
end entity audioInTest;

architecture rtl of audioInTest is
	component clocked_audio_input is
		generic (
			G_CAI_FIFO_DEPTH       : integer := 4;
			G_CAI_INCLUDE_CTRL_REG : integer := 0
		);
		port (
			reg_clk       : in  std_logic                     := 'X';             -- clk
			reg_reset     : in  std_logic                     := 'X';             -- reset
			aes_clk       : in  std_logic                     := 'X';             -- export
			aes_de        : in  std_logic                     := 'X';             -- export
			aes_ws        : in  std_logic                     := 'X';             -- export
			aes_data      : in  std_logic                     := 'X';             -- export
			aud_clk       : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			aud_ready     : in  std_logic                     := 'X';             -- ready
			aud_valid     : out std_logic;                                        -- valid
			aud_sop       : out std_logic;                                        -- startofpacket
			aud_eop       : out std_logic;                                        -- endofpacket
			aud_channel   : out std_logic_vector(7 downto 0);                     -- channel
			aud_data      : out std_logic_vector(23 downto 0);                    -- data
			channel0      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			channel1      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			fifo_status   : out std_logic_vector(7 downto 0);                     -- export
			fifo_reset    : in  std_logic                     := 'X';             -- export
			reg_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			reg_write     : in  std_logic                     := 'X';             -- write
			reg_writedata : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			reg_read      : in  std_logic                     := 'X';             -- read
			reg_readdata  : out std_logic_vector(7 downto 0)                      -- readdata
		);
	end component clocked_audio_input;

begin

	audiointest_inst : component clocked_audio_input
		generic map (
			G_CAI_FIFO_DEPTH       => 7,
			G_CAI_INCLUDE_CTRL_REG => 0
		)
		port map (
			reg_clk       => reg_clk,     --       control_clock.clk
			reg_reset     => reg_reset,   -- control_clock_reset.reset
			aes_clk       => aes_clk,     --   conduit_aes_audio.export
			aes_de        => aes_de,      --                    .export
			aes_ws        => aes_ws,      --                    .export
			aes_data      => aes_data,    --                    .export
			aud_clk       => aud_clk,     --          dout_clock.clk
			reset         => reset,       --    dout_clock_reset.reset
			aud_ready     => aud_ready,   --                dout.ready
			aud_valid     => aud_valid,   --                    .valid
			aud_sop       => aud_sop,     --                    .startofpacket
			aud_eop       => aud_eop,     --                    .endofpacket
			aud_channel   => aud_channel, --                    .channel
			aud_data      => aud_data,    --                    .data
			channel0      => channel0,    --     conduit_control.export
			channel1      => channel1,    --                    .export
			fifo_status   => fifo_status, --                    .export
			fifo_reset    => fifo_reset,  --                    .export
			reg_address   => "000",       --         (terminated)
			reg_write     => '0',         --         (terminated)
			reg_writedata => "00000000",  --         (terminated)
			reg_read      => '0',         --         (terminated)
			reg_readdata  => open         --         (terminated)
		);

end architecture rtl; -- of audioInTest
