-- megafunction wizard: %Clocked Audio Output Intel FPGA IP v20.1%
-- GENERATION: XML
-- outAudioTest.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity outAudioTest is
	port (
		reg_clk     : in  std_logic                     := '0';             --       control_clock.clk
		reg_reset   : in  std_logic                     := '0';             -- control_clock_reset.reset
		aud_clk     : in  std_logic                     := '0';             --           din_clock.clk
		reset       : in  std_logic                     := '0';             --     din_clock_reset.reset
		aud_ready   : out std_logic;                                        --                 din.ready
		aud_valid   : in  std_logic                     := '0';             --                    .valid
		aud_sop     : in  std_logic                     := '0';             --                    .startofpacket
		aud_eop     : in  std_logic                     := '0';             --                    .endofpacket
		aud_channel : in  std_logic_vector(7 downto 0)  := (others => '0'); --                    .channel
		aud_data    : in  std_logic_vector(23 downto 0) := (others => '0'); --                    .data
		aes_clk     : in  std_logic                     := '0';             --   conduit_aes_audio.export
		aes_de      : out std_logic;                                        --                    .export
		aes_ws      : out std_logic;                                        --                    .export
		aes_data    : out std_logic;                                        --                    .export
		channel0    : in  std_logic_vector(7 downto 0)  := (others => '0'); --     conduit_control.export
		channel1    : in  std_logic_vector(7 downto 0)  := (others => '0'); --                    .export
		fifo_status : out std_logic_vector(7 downto 0);                     --                    .export
		fifo_reset  : in  std_logic                     := '0'              --                    .export
	);
end entity outAudioTest;

architecture rtl of outAudioTest is
	component clocked_audio_output is
		generic (
			G_CAO_FIFO_DEPTH       : integer := 4;
			G_CAO_INCLUDE_CTRL_REG : integer := 0
		);
		port (
			reg_clk       : in  std_logic                     := 'X';             -- clk
			reg_reset     : in  std_logic                     := 'X';             -- reset
			aud_clk       : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			aud_ready     : out std_logic;                                        -- ready
			aud_valid     : in  std_logic                     := 'X';             -- valid
			aud_sop       : in  std_logic                     := 'X';             -- startofpacket
			aud_eop       : in  std_logic                     := 'X';             -- endofpacket
			aud_channel   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			aud_data      : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			aes_clk       : in  std_logic                     := 'X';             -- export
			aes_de        : out std_logic;                                        -- export
			aes_ws        : out std_logic;                                        -- export
			aes_data      : out std_logic;                                        -- export
			channel0      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			channel1      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			fifo_status   : out std_logic_vector(7 downto 0);                     -- export
			fifo_reset    : in  std_logic                     := 'X';             -- export
			reg_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			reg_write     : in  std_logic                     := 'X';             -- write
			reg_writedata : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			reg_read      : in  std_logic                     := 'X';             -- read
			reg_readdata  : out std_logic_vector(7 downto 0)                      -- readdata
		);
	end component clocked_audio_output;

begin

	outaudiotest_inst : component clocked_audio_output
		generic map (
			G_CAO_FIFO_DEPTH       => 7,
			G_CAO_INCLUDE_CTRL_REG => 0
		)
		port map (
			reg_clk       => reg_clk,     --       control_clock.clk
			reg_reset     => reg_reset,   -- control_clock_reset.reset
			aud_clk       => aud_clk,     --           din_clock.clk
			reset         => reset,       --     din_clock_reset.reset
			aud_ready     => aud_ready,   --                 din.ready
			aud_valid     => aud_valid,   --                    .valid
			aud_sop       => aud_sop,     --                    .startofpacket
			aud_eop       => aud_eop,     --                    .endofpacket
			aud_channel   => aud_channel, --                    .channel
			aud_data      => aud_data,    --                    .data
			aes_clk       => aes_clk,     --   conduit_aes_audio.export
			aes_de        => aes_de,      --                    .export
			aes_ws        => aes_ws,      --                    .export
			aes_data      => aes_data,    --                    .export
			channel0      => channel0,    --     conduit_control.export
			channel1      => channel1,    --                    .export
			fifo_status   => fifo_status, --                    .export
			fifo_reset    => fifo_reset,  --                    .export
			reg_address   => "000",       --         (terminated)
			reg_write     => '0',         --         (terminated)
			reg_writedata => "00000000",  --         (terminated)
			reg_read      => '0',         --         (terminated)
			reg_readdata  => open         --         (terminated)
		);

end architecture rtl; -- of outAudioTest
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2021 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="clocked_audio_output" version="20.1" >
-- Retrieval info: 	<generic name="FAMILY" value="Cyclone V" />
-- Retrieval info: 	<generic name="G_CAO_FIFO_DEPTH" value="7" />
-- Retrieval info: 	<generic name="G_CAO_INCLUDE_CTRL_REG" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : outAudioTest.vho
-- RELATED_FILES: outAudioTest.vhd, cao_fifo.v, cao_merge.v, cao_avalon.v, cao_registers.v, altera_cao_reset_synchronizer.v, clocked_audio_output.v
